module find_1_first(I,position,flag);
      input       [24:0]I;
      output	flag;
      output	[4:0]position;
      
      assign	flag=~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]
                      &~I[16]&~I[15]&~I[14]&~I[13]&~I[12]&~I[11]&~I[10]&~I[9]
      		    &~I[8]&~I[7]&~I[6]&~I[5]&~I[4]&~I[3]&~I[2]&~I[1]&~I[0];

      assign 	position[0]=(~I[24]&I[23])
                              |(~I[24]&~I[22]&I[21])
                              |(~I[24]&~I[22]&~I[20]&I[19])
      	                  |(~I[24]&~I[22]&~I[20]&~I[18]&I[17])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&I[15])
                               |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&I[13])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&I[11])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&I[9])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&~I[8]&I[7])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&~I[8]&~I[6]&I[5])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&~I[8]&~I[6]&~I[4]&I[3])
                              |(~I[24]&~I[22]&~I[20]&~I[18]&~I[16]&~I[14]&~I[12]&~I[10]&~I[8]&~I[6]&~I[4]&~I[2]&I[1]);

      assign	position[1]=(~I[24]&~I[23]&I[22])
                              |(~I[24]&~I[23]&I[21])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&I[18])
                              |(~I[24]&~I[23]&~I[20]&~I[19]&I[17])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&I[14])
                              |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&I[13])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&I[10])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&I[9])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&~I[8]&~I[7]&I[6])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&~I[8]&~I[7]&I[5])
                              |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&~I[8]&~I[7]&~I[4]&~I[3]&I[2])
      	                  |(~I[24]&~I[23]&~I[20]&~I[19]&~I[16]&~I[15]&~I[12]&~I[11]&~I[8]&~I[7]&~I[4]&~I[3]&I[1]);

      assign	position[2]=(~I[24]&~I[23]&~I[22]&~I[21]&I[20])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&I[19])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&I[18])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&I[17])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&I[12])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&I[11])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&I[10])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&I[9])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&~I[8]&~I[7]&~I[6]&~I[5]&I[4])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&~I[8]&~I[7]&~I[6]&~I[5]&I[3])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&~I[8]&~I[7]&~I[6]&~I[5]&I[2]) 
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[16]&~I[15]&~I[14]&~I[13]&~I[8]&~I[7]&~I[6]&~I[5]&I[1]);

      assign	position[3]=(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[16])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[15])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[14])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[13])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[12])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[11])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[10])
                              |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&I[9])
      	                  |(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&~I[8]&~I[7]&~I[6]&~I[5]&~I[4]&~I[3]&~I[2]&~I[1]&I[0]);

      assign	position[4]=(~I[24]&~I[23]&~I[22]&~I[21]&~I[20]&~I[19]&~I[18]&~I[17]&~I[16]&~I[15]
                        &~I[14]&~I[13]&~I[12]&~I[11]&~I[10]&~I[9])&(I[8]|I[7]|I[6]|I[5]|I[4]|I[3]|I[2]|I[1]|I[0]);

endmodule
